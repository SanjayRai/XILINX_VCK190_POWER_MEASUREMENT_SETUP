//Uncomment for NULL_BITSTREAM_DESIGN
//`define NULL_BITSTREAM_DESIGN
//`define SIMULATION_ONLY
